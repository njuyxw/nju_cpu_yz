module alu(
  input [3:0]ALUOP,
  input [31:0]inA,
  input [31:0]inB,
  output reg [31:0]aluout
  output reg zero,
  output reg overflow
);

  
endmodule 
